class operation;
  
  rand logic  a;
  rand logic  b;
  rand logic c;
  bit  sum;
  bit carry;
  
endclass
