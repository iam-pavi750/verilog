interface interfaces;
  
  logic d;
  logic clk;
  logic rst;
  bit q;
  
 endinterface
