class operation;
  
  logic  a;
 logic  b;
 logic c;
  bit  sum;
  bit carry;
  
endclass
