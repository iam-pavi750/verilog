class transaction;
  rand logic d;
   //logic clk;
   //logic rst;
  bit q;
endclass
